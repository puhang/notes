*---------- DMHT6016LFJ Spice Model ----------
.SUBCKT DMHT6016LFJ 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 NMOS L = 1E-006 W = 1E-006 
RD 10 1 0.006728 
RS 30 3 0.001 
RG 20 2 1.35 
CGS 2 3 8.475E-010 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 6E-010 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 5.378E+005 ETA = 0.001 VTO = 2.61 
+ TOX = 6E-008 NSUB = 1E+016 KP = 37.72 U0 = 400 KAPPA = 10 
.MODEL DCGD D CJO = 3.945E-010 VJ = 0.8 M = 0.6507 
.MODEL DSUB D IS = 2.448E-010 N = 1.248 RS = 0.006471 BV = 60 CJO = 5.274E-010 VJ = 0.8 M = 0.6 TT=2.2E-010
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMHT6016LFJ Spice Model v1.0 Last Revised 2016/11/23
